module MUX8to1(
    input [7:0] I,
    input [2:0] s,
    output [0:0] Y
    );
    assign Y = s[2]? (s[1]? (s[0]? I[7]:I[6]) : (s[0]? I[5]:I[4]))
                : (s[1]? (s[0]? I[3]:I[2]) : (s[0]? I[1]:I[0]));
endmodule



__________________________________________________________________________________________________________________________________________




module Mux8to1_tb ();

    reg [7:0] I;
    reg [2:0] s;
    wire Y;
    
    Mux8to1 uut (.I(I), .s(s), .Y(Y));
        initial begin
            
            I[7] = 0; I[6] = 0; I[5] = 0; I[4] = 0; I[3] = 0; I[2] = 0; I[1] = 0; I[0] = 1; s[2] = 0; s[1] = 0; s[0] = 0;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 1; I[4] = 1; I[3] = 1; I[2] = 1; I[1] = 1; I[0] = 0; s[2] = 0; s[1] = 0; s[0] = 0;
            #50;
            
            I[7] = 0; I[6] = 0; I[5] = 0; I[4] = 0; I[3] = 0; I[2] = 0; I[1] = 1; I[0] = 0; s[2] = 0; s[1] = 0; s[0] = 1;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 1; I[4] = 1; I[3] = 1; I[2] = 1; I[1] = 0; I[0] = 1; s[2] = 0; s[1] = 0; s[0] = 1;
            #50;
            
            I[7] = 0; I[6] = 0; I[5] = 0; I[4] = 0; I[3] = 0; I[2] = 1; I[1] = 0; I[0] = 0; s[2] = 0; s[1] = 1; s[0] = 0;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 1; I[4] = 1; I[3] = 1; I[2] = 0; I[1] = 1; I[0] = 1; s[2] = 0; s[1] = 1; s[0] = 0;
            #50;
            
            I[7] = 0; I[6] = 0; I[5] = 0; I[4] = 0; I[3] = 1; I[2] = 0; I[1] = 0; I[0] = 0; s[2] = 0; s[1] = 1; s[0] = 1;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 1; I[4] = 1; I[3] = 0; I[2] = 1; I[1] = 1; I[0] = 1; s[2] = 0; s[1] = 1; s[0] = 1;
            #50;
            
            I[7] = 0; I[6] = 0; I[5] = 0; I[4] = 1; I[3] = 0; I[2] = 0; I[1] = 0; I[0] = 0; s[2] = 1; s[1] = 0; s[0] = 0;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 1; I[4] = 0; I[3] = 1; I[2] = 1; I[1] = 1; I[0] = 1; s[2] = 1; s[1] = 0; s[0] = 0;
            #50;
            
            I[7] = 0; I[6] = 0; I[5] = 1; I[4] = 0; I[3] = 0; I[2] = 0; I[1] = 0; I[0] = 0; s[2] = 1; s[1] = 0; s[0] = 1;
            #50;
            I[7] = 1; I[6] = 1; I[5] = 0; I[4] = 1; I[3] = 1; I[2] = 1; I[1] = 1; I[0] = 1; s[2] = 1; s[1] = 0; s[0] = 1;
            #50;
            
            I[7] = 0; I[6] = 1; I[5] = 0; I[4] = 0; I[3] = 0; I[2] = 0; I[1] = 0; I[0] = 0; s[2] = 1; s[1] = 1; s[0] = 0;
            #50;
            I[7] = 1; I[6] = 0; I[5] = 1; I[4] = 1; I[3] = 1; I[2] = 1; I[1] = 1; I[0] = 1; s[2] = 1; s[1] = 1; s[0] = 0;
            #50;
            
            I[7] = 1; I[6] = 0; I[5] = 0; I[4] = 0; I[3] = 0; I[2] = 0; I[1] = 0; I[0] = 0; s[2] = 1; s[1] = 1; s[0] = 1;
            #50;
            I[7] = 0; I[6] = 1; I[5] = 1; I[4] = 1; I[3] = 1; I[2] = 1; I[1] = 1; I[0] = 1; s[2] = 1; s[1] = 1; s[0] = 1;
            #50;
        end
endmodule
